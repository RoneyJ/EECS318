

--test for CSA
entity testp4 is
end testp4;
