//receive logic module for the SSP of HW 3
//Josh Roney (jpr87)
module receive(
	input clear_b, pclk, sspclkin, sspfssin, ssprxd,
	output [7:0] rxdata,
	output sspoe_b, ssptxd, sspfssout, sspclkout
	);
endmodule;