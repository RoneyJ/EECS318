library verilog;
use verilog.vl_types.all;
entity Test_signed is
end Test_signed;
