--Structural FSM for HW4
--Josh Roney (jpr87)

entity structuralFSM is
	port(e,w,clock : in bit;
	     output : out bit);
end structuralFSM;
