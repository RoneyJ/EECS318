

--D Flip Flop for use by FSM
entity dff is
	port(d,clk : in bit;
	     q : out bit);
end DFF;
