library verilog;
use verilog.vl_types.all;
entity Add_9 is
    port(
        in1             : in     vl_logic_vector(8 downto 0);
        in2             : in     vl_logic_vector(8 downto 0);
        \out\           : out    vl_logic_vector(8 downto 0)
    );
end Add_9;
