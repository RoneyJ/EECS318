library verilog;
use verilog.vl_types.all;
entity P2_processor is
end P2_processor;
