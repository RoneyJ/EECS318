library verilog;
use verilog.vl_types.all;
entity Test_4x4 is
end Test_4x4;
