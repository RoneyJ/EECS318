library verilog;
use verilog.vl_types.all;
entity FSM_behav_test is
end FSM_behav_test;
