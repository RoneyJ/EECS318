library verilog;
use verilog.vl_types.all;
entity P1_processor is
end P1_processor;
