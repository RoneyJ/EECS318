library verilog;
use verilog.vl_types.all;
entity Test_shift_add is
end Test_shift_add;
