library verilog;
use verilog.vl_types.all;
entity \NOT\ is
    port(
        \out\           : out    vl_logic;
        \in\            : in     vl_logic
    );
end \NOT\;
