library verilog;
use verilog.vl_types.all;
entity ssp_test2 is
end ssp_test2;
