

--testbench for FSM
entity testP5b is
end testP5b;
