library verilog;
use verilog.vl_types.all;
entity Test_CSA is
end Test_CSA;
