

--test bench
entity testp2 is
end testp2;
