

--testbench for multiplier
entity testP1 is
end testP1;
