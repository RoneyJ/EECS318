--Behavioral FSM for HW4
--Josh Roney (jpr87)
entity behavioralFSM is
	port(e,w,clk : in bit;
	     o : out bit);
end entity;
