library verilog;
use verilog.vl_types.all;
entity ssp_test1 is
end ssp_test1;
