 


--full adder for use of multiplier
entity fa is
	port(a,b,cin : in bit;
	     cout,s : out bit);
end entity;
