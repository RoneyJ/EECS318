library verilog;
use verilog.vl_types.all;
entity FSM_Struc_Test is
end FSM_Struc_Test;
