library verilog;
use verilog.vl_types.all;
entity testHandshake is
end testHandshake;
