library verilog;
use verilog.vl_types.all;
entity Test_adder is
end Test_adder;
