library verilog;
use verilog.vl_types.all;
entity testFreeCell is
end testFreeCell;
