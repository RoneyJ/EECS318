library verilog;
use verilog.vl_types.all;
entity P3_processor is
end P3_processor;
