

--test bench
entity testp3 is
end testp3;
