

--testbench for FSM
entity testP5s is
end testP5s;
