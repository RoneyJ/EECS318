library verilog;
use verilog.vl_types.all;
entity test_tfifo is
end test_tfifo;
